
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity HAZARD_DETECTION_UNIT is
PORT(a:IN STD_LOGIC
);
end HAZARD_DETECTION_UNIT;

architecture Behavioral of HAZARD_DETECTION_UNIT is

begin


end Behavioral;

