library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity program_counter is
port(pc_in: in std_logic_vector(15 downto 0);
pc_out: out std_logic_vector(15 downto 0);

end program_counter;

architecture Behavioral of program_counter is

begin


end Behavioral;

