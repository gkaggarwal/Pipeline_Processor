
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity CONTROLLER is
PORT(A: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
OUTPUT: OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
);
end CONTROLLER;

architecture Behavioral of CONTROLLER is
begin
PROCESS(A)
BEGIN
IF (A(15 DOWNTO 12)="0000" AND A(1 DOWNTO 0)="00" )THEN
OUTPUT(5 DOWNTO 0)<="000001";
OUTPUT(11 DOWNTO 6)<="100000";
OUTPUT(17 DOWNTO 12)<="000000";
OUTPUT(23 DOWNTO 18)<="000001";
ELSIF((A(15 DOWNTO 12)="0000"  OR A(15 DOWNTO 12)="0010") AND A(1 DOWNTO 0)="01")THEN
OUTPUT(5 DOWNTO 0)<="000001";
OUTPUT(11 DOWNTO 6)<="100000";
OUTPUT(17 DOWNTO 12)<="000000";
OUTPUT(23 DOWNTO 18)<="000011";
ELSIF((A(15 DOWNTO 12)="0000" OR A(15 DOWNTO 12)="0010") AND A(1 DOWNTO 0)="10")THEN
OUTPUT(5 DOWNTO 0)<="000001";
OUTPUT(11 DOWNTO 6)<="100000";
OUTPUT(17 DOWNTO 12)<="000000";
OUTPUT(23 DOWNTO 18)<="000101";
ELSIF(A(15 DOWNTO 12)="0001" OR A(15 DOWNTO 12)="0010")THEN
OUTPUT(5 DOWNTO 0)<="000001";
OUTPUT(11 DOWNTO 6)<="100000";
OUTPUT(17 DOWNTO 12)<="000000";
OUTPUT(23 DOWNTO 18)<="000001";
ELSIF(A(15 DOWNTO 12)="0011")THEN
OUTPUT(5 DOWNTO 0)<="000000";
OUTPUT(11 DOWNTO 6)<="100000";
OUTPUT(17 DOWNTO 12)<="000000";
OUTPUT(23 DOWNTO 18)<="000001";
ELSIF(A(15 DOWNTO 12)="0100")THEN
OUTPUT(5 DOWNTO 0)<="000001";
OUTPUT(11 DOWNTO 6)<="100000";
OUTPUT(17 DOWNTO 12)<="000010";
OUTPUT(23 DOWNTO 18)<="001001";
ELSIF(A(15 DOWNTO 12)="0101")THEN
OUTPUT(5 DOWNTO 0)<="000011";
OUTPUT(11 DOWNTO 6)<="100000";
OUTPUT(17 DOWNTO 12)<="000001";
OUTPUT(23 DOWNTO 18)<="000000";
ELSIF(A(15 DOWNTO 12)="1100")THEN
OUTPUT(5 DOWNTO 0)<="000011";
OUTPUT(11 DOWNTO 6)<="100000";
OUTPUT(17 DOWNTO 12)<="000101";
OUTPUT(23 DOWNTO 18)<="000000";
ELSIF(A(15 DOWNTO 12)="1000")THEN
OUTPUT(5 DOWNTO 0)<="000000";
OUTPUT(11 DOWNTO 6)<="100001";
OUTPUT(17 DOWNTO 12)<="000000";
OUTPUT(23 DOWNTO 18)<="010001";
ELSIF(A(15 DOWNTO 12)="1001")THEN
OUTPUT(5 DOWNTO 0)<="000001";
OUTPUT(11 DOWNTO 6)<="100010";
OUTPUT(17 DOWNTO 12)<="000000";
OUTPUT(23 DOWNTO 18)<="010001";
ELSIF(A(15 DOWNTO 12)="0110")THEN
OUTPUT(5 DOWNTO 0)<="000011";
OUTPUT(11 DOWNTO 6)<="010100";
OUTPUT(17 DOWNTO 12)<="000010";
OUTPUT(23 DOWNTO 18)<="101001";
ELSIF(A(15 DOWNTO 12)="0111")THEN
OUTPUT(5 DOWNTO 0)<="000111";
OUTPUT(11 DOWNTO 6)<="010100";
OUTPUT(17 DOWNTO 12)<="001001";
OUTPUT(23 DOWNTO 18)<="000000";
ELSE
OUTPUT(5 DOWNTO 0)<="000000";
OUTPUT(11 DOWNTO 6)<="100000";
OUTPUT(17 DOWNTO 12)<="000000";
OUTPUT(23 DOWNTO 18)<="000000";
END IF;
END PROCESS;
end Behavioral;

